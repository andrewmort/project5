library verilog;
use verilog.vl_types.all;
entity bsr_tb is
end bsr_tb;
