library verilog;
use verilog.vl_types.all;
entity s9234 is
    port(
        CK              : in     vl_logic;
        g89             : in     vl_logic;
        g94             : in     vl_logic;
        g98             : in     vl_logic;
        g102            : in     vl_logic;
        g107            : in     vl_logic;
        g301            : in     vl_logic;
        g306            : in     vl_logic;
        g310            : in     vl_logic;
        g314            : in     vl_logic;
        g319            : in     vl_logic;
        g557            : in     vl_logic;
        g558            : in     vl_logic;
        g559            : in     vl_logic;
        g560            : in     vl_logic;
        g561            : in     vl_logic;
        g562            : in     vl_logic;
        g563            : in     vl_logic;
        g564            : in     vl_logic;
        g705            : in     vl_logic;
        g639            : in     vl_logic;
        g567            : in     vl_logic;
        g45             : in     vl_logic;
        g42             : in     vl_logic;
        g39             : in     vl_logic;
        g702            : in     vl_logic;
        g32             : in     vl_logic;
        g38             : in     vl_logic;
        g46             : in     vl_logic;
        g36             : in     vl_logic;
        g47             : in     vl_logic;
        g40             : in     vl_logic;
        g37             : in     vl_logic;
        g41             : in     vl_logic;
        g22             : in     vl_logic;
        g44             : in     vl_logic;
        g23             : in     vl_logic;
        g2584           : out    vl_logic;
        g3222           : out    vl_logic;
        g3600           : out    vl_logic;
        g4307           : out    vl_logic;
        g4321           : out    vl_logic;
        g4422           : out    vl_logic;
        g4809           : out    vl_logic;
        g5137           : out    vl_logic;
        g5468           : out    vl_logic;
        g5469           : out    vl_logic;
        g5692           : out    vl_logic;
        g6282           : out    vl_logic;
        g6284           : out    vl_logic;
        g6360           : out    vl_logic;
        g6362           : out    vl_logic;
        g6364           : out    vl_logic;
        g6366           : out    vl_logic;
        g6368           : out    vl_logic;
        g6370           : out    vl_logic;
        g6372           : out    vl_logic;
        g6374           : out    vl_logic;
        g6728           : out    vl_logic;
        g1290           : out    vl_logic;
        g4121           : out    vl_logic;
        g4108           : out    vl_logic;
        g4106           : out    vl_logic;
        g4103           : out    vl_logic;
        g1293           : out    vl_logic;
        g4099           : out    vl_logic;
        g4102           : out    vl_logic;
        g4109           : out    vl_logic;
        g4100           : out    vl_logic;
        g4112           : out    vl_logic;
        g4105           : out    vl_logic;
        g4101           : out    vl_logic;
        g4110           : out    vl_logic;
        g4104           : out    vl_logic;
        g4107           : out    vl_logic;
        g4098           : out    vl_logic
    );
end s9234;
