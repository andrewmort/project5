library verilog;
use verilog.vl_types.all;
entity TB_modulename is
end TB_modulename;
