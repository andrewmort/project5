library verilog;
use verilog.vl_types.all;
entity udff_r is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end udff_r;
