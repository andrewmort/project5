library verilog;
use verilog.vl_types.all;
entity s9234_tap is
    port(
        TDO             : out    vl_logic;
        CK              : in     vl_logic;
        TDI             : in     vl_logic;
        TMS             : in     vl_logic;
        TRST_b          : in     vl_logic;
        g89i            : in     vl_logic;
        g94i            : in     vl_logic;
        g98i            : in     vl_logic;
        g102i           : in     vl_logic;
        g107i           : in     vl_logic;
        g301i           : in     vl_logic;
        g306i           : in     vl_logic;
        g310i           : in     vl_logic;
        g314i           : in     vl_logic;
        g319i           : in     vl_logic;
        g557i           : in     vl_logic;
        g558i           : in     vl_logic;
        g559i           : in     vl_logic;
        g560i           : in     vl_logic;
        g561i           : in     vl_logic;
        g562i           : in     vl_logic;
        g563i           : in     vl_logic;
        g564i           : in     vl_logic;
        g705i           : in     vl_logic;
        g639i           : in     vl_logic;
        g567i           : in     vl_logic;
        g45i            : in     vl_logic;
        g42i            : in     vl_logic;
        g39i            : in     vl_logic;
        g702i           : in     vl_logic;
        g32i            : in     vl_logic;
        g38i            : in     vl_logic;
        g46i            : in     vl_logic;
        g36i            : in     vl_logic;
        g47i            : in     vl_logic;
        g40i            : in     vl_logic;
        g37i            : in     vl_logic;
        g41i            : in     vl_logic;
        g22i            : in     vl_logic;
        g44i            : in     vl_logic;
        g23i            : in     vl_logic;
        g2584           : out    vl_logic;
        g3222           : out    vl_logic;
        g3600           : out    vl_logic;
        g4307           : out    vl_logic;
        g4321           : out    vl_logic;
        g4422           : out    vl_logic;
        g4809           : out    vl_logic;
        g5137           : out    vl_logic;
        g5468           : out    vl_logic;
        g5469           : out    vl_logic;
        g5692           : out    vl_logic;
        g6282           : out    vl_logic;
        g6284           : out    vl_logic;
        g6360           : out    vl_logic;
        g6362           : out    vl_logic;
        g6364           : out    vl_logic;
        g6366           : out    vl_logic;
        g6368           : out    vl_logic;
        g6370           : out    vl_logic;
        g6372           : out    vl_logic;
        g6374           : out    vl_logic;
        g6728           : out    vl_logic;
        g1290           : out    vl_logic;
        g4121           : out    vl_logic;
        g4108           : out    vl_logic;
        g4106           : out    vl_logic;
        g4103           : out    vl_logic;
        g1293           : out    vl_logic;
        g4099           : out    vl_logic;
        g4102           : out    vl_logic;
        g4109           : out    vl_logic;
        g4100           : out    vl_logic;
        g4112           : out    vl_logic;
        g4105           : out    vl_logic;
        g4101           : out    vl_logic;
        g4110           : out    vl_logic;
        g4104           : out    vl_logic;
        g4107           : out    vl_logic;
        g4098           : out    vl_logic
    );
end s9234_tap;
