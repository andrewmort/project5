library verilog;
use verilog.vl_types.all;
entity normaltb is
end normaltb;
